-- Copyright (C) 2020  Intel Corporation. All rights reserved.
-- Your use of Intel Corporation's design tools, logic functions 
-- and other software and tools, and any partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Intel Program License 
-- Subscription Agreement, the Intel Quartus Prime License Agreement,
-- the Intel FPGA IP License Agreement, or other applicable license
-- agreement, including, without limitation, that your use is for
-- the sole purpose of programming logic devices manufactured by
-- Intel and sold by Intel or its authorized distributors.  Please
-- refer to the applicable agreement for further details, at
-- https://fpgasoftware.intel.com/eula.

-- PROGRAM		"Quartus Prime"
-- VERSION		"Version 20.1.1 Build 720 11/11/2020 SJ Lite Edition"
-- CREATED		"Fri Oct 27 12:26:59 2023"

LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY Synth IS 
	PORT
	(
		clk :  IN  STD_LOGIC;
		D :  IN  STD_LOGIC;
		E :  IN  STD_LOGIC;
		F :  IN  STD_LOGIC;
		G :  IN  STD_LOGIC;
		A :  IN  STD_LOGIC;
		speed_up :  IN  STD_LOGIC;
		nrst :  IN  STD_LOGIC;
		C :  IN  STD_LOGIC;
		en :  IN  STD_LOGIC_VECTOR(1 DOWNTO 0);
		sequence_enab :  IN  STD_LOGIC_VECTOR(1 DOWNTO 0);
		i_data :  OUT  STD_LOGIC_VECTOR(8 DOWNTO 0);
		seg6 :  OUT  STD_LOGIC;
		seg5 :  OUT  STD_LOGIC;
		seg4 :  OUT  STD_LOGIC;
		seg3 :  OUT  STD_LOGIC;
		seg2 :  OUT  STD_LOGIC;
		seg1 :  OUT  STD_LOGIC;
		seg0 :  OUT  STD_LOGIC;
		seg16 :  OUT  STD_LOGIC;
		seg15 :  OUT  STD_LOGIC;
		seg14 :  OUT  STD_LOGIC;
		seg13 :  OUT  STD_LOGIC;
		seg12 :  OUT  STD_LOGIC;
		seg11 :  OUT  STD_LOGIC;
		seg10 :  OUT  STD_LOGIC
	);
END Synth;

ARCHITECTURE bdf_type OF Synth IS 

COMPONENT monothonic_synth
	PORT(C : IN STD_LOGIC;
		 D : IN STD_LOGIC;
		 E : IN STD_LOGIC;
		 F : IN STD_LOGIC;
		 G : IN STD_LOGIC;
		 A : IN STD_LOGIC;
		 nrst : IN STD_LOGIC;
		 clk : IN STD_LOGIC;
		 speed_up : IN STD_LOGIC;
		 en : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
		 sequence_enab : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
		 BPM_dis : OUT STD_LOGIC_VECTOR(8 DOWNTO 0);
		 i_data : OUT STD_LOGIC_VECTOR(8 DOWNTO 0)
	);
END COMPONENT;

COMPONENT toseg
	PORT(bcd : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		 seg : OUT STD_LOGIC_VECTOR(6 DOWNTO 0)
	);
END COMPONENT;

SIGNAL	BPM_dis :  STD_LOGIC_VECTOR(8 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_12 :  STD_LOGIC_VECTOR(6 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_13 :  STD_LOGIC_VECTOR(6 DOWNTO 0);


BEGIN 
seg6 <= SYNTHESIZED_WIRE_12(6);
seg5 <= SYNTHESIZED_WIRE_12(5);
seg4 <= SYNTHESIZED_WIRE_12(4);
seg3 <= SYNTHESIZED_WIRE_12(3);
seg2 <= SYNTHESIZED_WIRE_12(2);
seg1 <= SYNTHESIZED_WIRE_12(1);
seg0 <= SYNTHESIZED_WIRE_12(0);
seg16 <= SYNTHESIZED_WIRE_13(6);
seg15 <= SYNTHESIZED_WIRE_13(5);
seg14 <= SYNTHESIZED_WIRE_13(4);
seg13 <= SYNTHESIZED_WIRE_13(3);
seg12 <= SYNTHESIZED_WIRE_13(2);
seg11 <= SYNTHESIZED_WIRE_13(1);
seg10 <= SYNTHESIZED_WIRE_13(0);



b2v_inst : monothonic_synth
PORT MAP(C => C,
		 D => D,
		 E => E,
		 F => F,
		 G => G,
		 A => A,
		 nrst => nrst,
		 clk => clk,
		 speed_up => speed_up,
		 en => en,
		 sequence_enab => sequence_enab,
		 BPM_dis => BPM_dis,
		 i_data => i_data);


b2v_inst1 : toseg
PORT MAP(bcd => BPM_dis(3 DOWNTO 0),
		 seg => SYNTHESIZED_WIRE_12);


b2v_inst2 : toseg
PORT MAP(bcd => BPM_dis(7 DOWNTO 4),
		 seg => SYNTHESIZED_WIRE_13);



BPM_dis(8) <= '0';
END bdf_type;